../../jtag_reset.vhd