-- shamt_roms.vhd
-- Copyright (C) 2015 VectorBlox Computing, Inc.

-- synthesis library vbx_lib
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;
use work.util_pkg.all;
use work.isa_pkg.all;
use work.architecture_pkg.all;
use work.component_pkg.all;

entity byte_shamt_rom is
  port
    (
      shamt_trunc        : in  std_logic_vector(2 downto 0);
      shiftl             : in  std_logic;
      byte_shamt_rom_out : out std_logic_vector(8 downto 0)
      );
end byte_shamt_rom;

architecture syn of byte_shamt_rom is
  signal shiftl_shamt : std_logic_vector(3 downto 0);
begin

  shiftl_shamt <= shiftl & shamt_trunc;
  with shiftl_shamt select
    byte_shamt_rom_out(8 downto 0) <=
    "100000000" when "0000",
    "010000000" when "0001",
    "001000000" when "0010",
    "000100000" when "0011",
    "000010000" when "0100",
    "000001000" when "0101",
    "000000100" when "0110",
    "000000010" when "0111",
    "000000001" when "1000",
    "000000010" when "1001",
    "000000100" when "1010",
    "000001000" when "1011",
    "000010000" when "1100",
    "000100000" when "1101",
    "001000000" when "1110",
    "010000000" when "1111",
    "000000000" when others;
  
end syn;


-- synthesis library vbx_lib
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;
use work.util_pkg.all;
use work.isa_pkg.all;
use work.architecture_pkg.all;
use work.component_pkg.all;

entity half_shamt_rom is
  port
    (
      shamt_trunc        : in  std_logic_vector(3 downto 0);
      shiftl             : in  std_logic;
      half_shamt_rom_out : out std_logic_vector(17 downto 0)
      );
end half_shamt_rom;

architecture syn of half_shamt_rom is
  signal shiftl_shamt : std_logic_vector(4 downto 0);
begin
  half_shamt_rom_out(17) <= '0';

  shiftl_shamt <= shiftl & shamt_trunc;
  with shiftl_shamt select
    half_shamt_rom_out(16 downto 0) <=
    "10000000000000000" when "00000",
    "01000000000000000" when "00001",
    "00100000000000000" when "00010",
    "00010000000000000" when "00011",
    "00001000000000000" when "00100",
    "00000100000000000" when "00101",
    "00000010000000000" when "00110",
    "00000001000000000" when "00111",
    "00000000100000000" when "01000",
    "00000000010000000" when "01001",
    "00000000001000000" when "01010",
    "00000000000100000" when "01011",
    "00000000000010000" when "01100",
    "00000000000001000" when "01101",
    "00000000000000100" when "01110",
    "00000000000000010" when "01111",
    "00000000000000001" when "10000",
    "00000000000000010" when "10001",
    "00000000000000100" when "10010",
    "00000000000001000" when "10011",
    "00000000000010000" when "10100",
    "00000000000100000" when "10101",
    "00000000001000000" when "10110",
    "00000000010000000" when "10111",
    "00000000100000000" when "11000",
    "00000001000000000" when "11001",
    "00000010000000000" when "11010",
    "00000100000000000" when "11011",
    "00001000000000000" when "11100",
    "00010000000000000" when "11101",
    "00100000000000000" when "11110",
    "01000000000000000" when "11111",
    "00000000000000000" when others;
  
end syn;


-- synthesis library vbx_lib
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;
use work.util_pkg.all;
use work.isa_pkg.all;
use work.architecture_pkg.all;
use work.component_pkg.all;

entity word_shamt_rom is
  port
    (
      shamt_trunc        : in  std_logic_vector(4 downto 0);
      shiftl             : in  std_logic;
      word_shamt_rom_out : out std_logic_vector(33 downto 0)
      );
end word_shamt_rom;

architecture syn of word_shamt_rom is
  signal shiftl_shamt : std_logic_vector(5 downto 0);
begin
  word_shamt_rom_out(33) <= '0';

  shiftl_shamt <= shiftl & shamt_trunc;
  with shiftl_shamt select
    word_shamt_rom_out(32 downto 0) <=
    "100000000000000000000000000000000" when "000000",
    "010000000000000000000000000000000" when "000001",
    "001000000000000000000000000000000" when "000010",
    "000100000000000000000000000000000" when "000011",
    "000010000000000000000000000000000" when "000100",
    "000001000000000000000000000000000" when "000101",
    "000000100000000000000000000000000" when "000110",
    "000000010000000000000000000000000" when "000111",
    "000000001000000000000000000000000" when "001000",
    "000000000100000000000000000000000" when "001001",
    "000000000010000000000000000000000" when "001010",
    "000000000001000000000000000000000" when "001011",
    "000000000000100000000000000000000" when "001100",
    "000000000000010000000000000000000" when "001101",
    "000000000000001000000000000000000" when "001110",
    "000000000000000100000000000000000" when "001111",
    "000000000000000010000000000000000" when "010000",
    "000000000000000001000000000000000" when "010001",
    "000000000000000000100000000000000" when "010010",
    "000000000000000000010000000000000" when "010011",
    "000000000000000000001000000000000" when "010100",
    "000000000000000000000100000000000" when "010101",
    "000000000000000000000010000000000" when "010110",
    "000000000000000000000001000000000" when "010111",
    "000000000000000000000000100000000" when "011000",
    "000000000000000000000000010000000" when "011001",
    "000000000000000000000000001000000" when "011010",
    "000000000000000000000000000100000" when "011011",
    "000000000000000000000000000010000" when "011100",
    "000000000000000000000000000001000" when "011101",
    "000000000000000000000000000000100" when "011110",
    "000000000000000000000000000000010" when "011111",
    "000000000000000000000000000000001" when "100000",
    "000000000000000000000000000000010" when "100001",
    "000000000000000000000000000000100" when "100010",
    "000000000000000000000000000001000" when "100011",
    "000000000000000000000000000010000" when "100100",
    "000000000000000000000000000100000" when "100101",
    "000000000000000000000000001000000" when "100110",
    "000000000000000000000000010000000" when "100111",
    "000000000000000000000000100000000" when "101000",
    "000000000000000000000001000000000" when "101001",
    "000000000000000000000010000000000" when "101010",
    "000000000000000000000100000000000" when "101011",
    "000000000000000000001000000000000" when "101100",
    "000000000000000000010000000000000" when "101101",
    "000000000000000000100000000000000" when "101110",
    "000000000000000001000000000000000" when "101111",
    "000000000000000010000000000000000" when "110000",
    "000000000000000100000000000000000" when "110001",
    "000000000000001000000000000000000" when "110010",
    "000000000000010000000000000000000" when "110011",
    "000000000000100000000000000000000" when "110100",
    "000000000001000000000000000000000" when "110101",
    "000000000010000000000000000000000" when "110110",
    "000000000100000000000000000000000" when "110111",
    "000000001000000000000000000000000" when "111000",
    "000000010000000000000000000000000" when "111001",
    "000000100000000000000000000000000" when "111010",
    "000001000000000000000000000000000" when "111011",
    "000010000000000000000000000000000" when "111100",
    "000100000000000000000000000000000" when "111101",
    "001000000000000000000000000000000" when "111110",
    "010000000000000000000000000000000" when "111111",
    "000000000000000000000000000000000" when others;
  
end syn;
