../../../rtl/a4l_master.vhd