../../rtl/lve_ci.vhd