../../rtl/4port_mem.vhd