../../../rtl/a4l_instruction_master.vhd