../../iram_xilinx.vhd