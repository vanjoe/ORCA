../../rtl/apb_to_ram.vhd