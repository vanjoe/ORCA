../../rtl/axi_wrapper.vhd