../../../rtl/cache.vhd